// timmer,  generates one pulse of clk period width each PERIOD count of clk

// parameter 2^WIDTH must be bigger then PERIOD
// parameter PERIOD must be bigger then 2

module timer #(parameter WIDTH = 32, parameter PERIOD = 1000)(
	input  clk,
	output reg out
	);
	
// TASK 1a: here is a place for your code

endmodule